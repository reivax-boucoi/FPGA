module vga(
    input clk,
    input clear,
    input [7:0] sw
    );


endmodule
